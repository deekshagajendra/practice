
Checking git pull
