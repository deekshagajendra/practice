bejbvjk
